`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 23.05.2024 14:37:21
// Design Name: 
// Module Name: Four_wires
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Four_wires(input a,b,c, output w,x,y,z);
assign w=a;
assign x=b;
assign y=b;
assign z=c;

endmodule
